//`timescale 1ns/1ns
//
//module tb9;
//
//logic enter, clk, overflow, tab, rst;
//logic [1:0] state, nextstate;
//
//autoupd autoupd (.clk(clk), .addr()addr, .in(in), .out(out), .state(state), .nextstate(nextstate), .rst(rst));
//
//initial begin
// rst = 1;
// clk = 0;
//end
//
//
//endmodule