// just for info

module ascii ();

enum logic [7:0]
{
NULL=8'd0,
SOH=8'd1,
STX=8'd	2	,
ETX=8'd	3	,
EOT=8'd	4	,
ENQ=8'd	5	,
ACK=8'd	6	,
BEL=8'd	7	,
BS=8'd	8	,
HT=8'd	9	,
LF=8'd	10	,
VT=8'd	11	,
FF=8'd	12	,
CR=8'd	13	,
SO=8'd	14	,
SI=8'd	15	,
DLE=8'd	16	,
DC1=8'd	17	,
DC2=8'd	18	,
DC3=8'd	19	,
DC4=8'd	20	,
NAK=8'd	21	,
SYN=8'd	22	,
ETB=8'd	23	,
CAN=8'd	24	,
EM=8'd	25	,
SUB=8'd	26	,
ESC=8'd	27	,
FS=8'd	28	,
GS=8'd	29	,
RS=8'd	30	,
US=8'd	31	,
Space=8'd	32	,
Exclamation=8'd	33	,
quotes	=8'd	34	,
OCTOTHORPE	=8'd	35	,
dollar	=8'd	36	,
percent	=8'd	37	,
AMPERSAND	=8'd	38	,
APOSTROPHE	=8'd	39	,
OPENPARENTHESIS	=8'd	40	,
CLOSEPARENTHESIS	=8'd	41	,
ASTERISK	=8'd	42	,
PLUS	=8'd	43	,
COMMA	=8'd	44	,
MINUS	=8'd	45	,
DOT	=8'd	46	,
FORWARDSLASH	=8'd	47	,
zero	=8'd	48	,
one	=8'd	49	,
two	=8'd	50	,
three	=8'd	51	,
four	=8'd	52	,
five	=8'd	53	,
six	=8'd	54	,
seven	=8'd	55	,
eight	=8'd	56	,
nine	=8'd	57	,
COLON	=8'd	58	,
SEMICOLON	=8'd	59	,
LESS	=8'd	60	,
EQUALS	=8'd	61	,
GREATER	=8'd	62	,
QUESTION	=8'd	63	,
ATORAT	=8'd	64	,
A	=8'd	65	,
B	=8'd	66	,
C	=8'd	67	,
D	=8'd	68	,
E	=8'd	69	,
F	=8'd	70	,
G	=8'd	71	,
H	=8'd	72	,
I	=8'd	73	,
J	=8'd	74	,
K	=8'd	75	,
L	=8'd	76	,
M	=8'd	77	,
N	=8'd	78	,
O	=8'd	79	,
P	=8'd	80	,
Q	=8'd	81	,
R	=8'd	82	,
S	=8'd	83	,
T	=8'd	84	,
U	=8'd	85	,
V	=8'd	86	,
W	=8'd	87	,
X	=8'd	88	,
Y	=8'd	89	,
Z	=8'd	90	,
squareright	=8'd	91	,
backslash	=8'd	92	,
squareleft	=8'd	93	,
CARET	=8'd	94	,
UNDERSCORE	=8'd	95	,
ACUTE	=8'd	96	,
a	=8'd	97	,
b	=8'd	98	,
c	=8'd	99	,
d	=8'd	100	,
e	=8'd	101	,
f	=8'd	102	,
g	=8'd	103	,
h	=8'd	104	,
i	=8'd	105	,
j	=8'd	106	,
k	=8'd	107	,
l	=8'd	108	,
m	=8'd	109	,
n	=8'd	110	,
o	=8'd	111	,
p	=8'd	112	,
q	=8'd	113	,
r	=8'd	114	,
s	=8'd	115	,
t	=8'd	116	,
u	=8'd	117	,
v	=8'd	118	,
w	=8'd	119	,
x	=8'd	120	,
y	=8'd	121	,
z	=8'd	122	,
leftcurly	=8'd	123	,
VERTICALBAR	=8'd	124	,
rightcurly	=8'd	125	,
TILDE	=8'd	126	,
DEL	=8'd	127
} ascii;


endmodule